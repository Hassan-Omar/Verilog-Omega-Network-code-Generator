module OmegaNetwork(input [7:0] InDat, input CLK, output [7:0]  outData);
    wire WS0_0;
    wire WS0_1;
    wire WS0_2;
    wire WS0_3;
    wire WS0_4;
    wire WS0_5;
    wire WS0_6;
    wire WS0_7;
    wire WS1_0;
    wire WS1_1;
    wire WS1_2;
    wire WS1_3;
    wire WS1_4;
    wire WS1_5;
    wire WS1_6;
    wire WS1_7;
    wire WS2_0;
    wire WS2_1;
    wire WS2_2;
    wire WS2_3;
    wire WS2_4;
    wire WS2_5;
    wire WS2_6;
    wire WS2_7;
    Banyan2_2 ins_Banyn0_0(InDat[7], InDat[6], WS0_0, WS0_1, CLK);
    Banyan2_2 ins_Banyn1_0(InDat[5], InDat[4], WS0_2, WS0_3, CLK);
    Banyan2_2 ins_Banyn2_0(InDat[3], InDat[2], WS0_4, WS0_5, CLK);
    Banyan2_2 ins_Banyn3_0(InDat[1], InDat[0], WS0_6, WS0_7, CLK);
    Banyan2_2 ins_Banyn0_1(WS0_0, WS0_4, WS1_0, WS1_1, CLK);
    Banyan2_2 ins_Banyn1_1(WS0_1, WS0_5, WS1_2, WS1_3, CLK);
    Banyan2_2 ins_Banyn2_1(WS0_2, WS0_6, WS1_4, WS1_5, CLK);
    Banyan2_2 ins_Banyn3_1(WS0_3, WS0_7, WS1_6, WS1_7, CLK);
    Banyan2_2 ins_Banyn0_2(WS1_0, WS1_4, outData[7], outData[6], CLK);
    Banyan2_2 ins_Banyn1_2(WS1_1, WS1_5, outData[5], outData[4], CLK);
    Banyan2_2 ins_Banyn2_2(WS1_2, WS1_6, outData[3], outData[2], CLK);
    Banyan2_2 ins_Banyn3_2(WS1_3, WS1_7, outData[1], outData[0], CLK);
endmodule